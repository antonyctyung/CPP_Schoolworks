** Profile: "SCHEMATIC1-ece2200_sim_m1"  [ D:\Documents\workspace\CPP_Schoolworks\ECE2200\PSpiceActivity\ece2200_m1-PSpiceFiles\SCHEMATIC1\ece2200_sim_m1.sim ] 

** Creating circuit file "ece2200_sim_m1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ece2200_m1-pspicefiles/ece2200_m1.lib" 
* From [PSPICE NETLIST] section of C:\Users\Antony Yung\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 .1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

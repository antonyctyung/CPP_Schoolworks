** Profile: "SCHEMATIC1-sim"  [ D:\Documents\workspace\CPP_Schoolworks\ECE2200L\ECE2200L_Lab3\ECE2200L_Lab3_PSpice\ece2200l_lab3-pspicefiles\schematic1\sim.sim ] 

** Creating circuit file "sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Antony Yung\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC LIN 1 60 60
.STEP LIN PARAM vin -100 100 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

ECE2101L Lab7 Part B2: Measuring OUTPUT impedance of a black box with 130 Ohm resistor
* Author: Choi Tim Antony Yung
* Simulation using 130ohm resistor

.INCLUDE blackbox.cir

XBOX v0 0 BOX
R0 v0 0 130
.AC LIN 1 60 60
.PRINT AC v(v0)

.END
